Photodiode
.include lm324.txt
CJ 1 0 11p
C1 1 4 3.3p
C2 2 0 1u
r1 1 4 1.4Meg
r2 2 3 13.7k
r3 2 0 280
x1 2 1 3 0 4 LM324
vcc 3 0 +5
vref 2 0 0.1
I1 1 0 dc 1.5u ac 1
.ac dec 10 10 100Meg
.control
run
plot vdb(4)
.endc
.end

