Schmitt Trigger
.include ua741.txt
.SUBCKT ZENER_12 1 2 
D1 1 2 DF 
DZ 3 1 DR 
VZ 2 3 3.5
.MODEL DF D ( IS=27.5p 
+RS=0.620
+N=1.10
+CJO=78.3p
+VJ=1.00
+M=0.330 
+TT=50.1n) 
.MODEL DR D ( IS=5.49f RS=50 N=1.77 ) 
.ends
X1 1 2 3 4 5 ua741
vcc 3 0 +15v
vdd 4 0 -15v
r1 5 6 1k
r2 6 1 10k
r3 1 8 10k
x2 6 7 ZENER_12 
x3 0 7 ZENER_12
va 8 0 3v
*voltage input 
vin 2 0 sin(0 6v 1k 0 0)
.tran 0.001ms 10ms
.control
run
plot v(6)
plot v(6) vs v(2)
.endc
.end